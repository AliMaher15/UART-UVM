interface uart_rx_system_if (input clk);

    bit    res_n;    //output
    
endinterface : uart_rx_system_if
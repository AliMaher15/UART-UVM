package uart_rx_seq_pkg ;
    
	import uvm_pkg::*;
	`include "uvm_macros.svh"

    import uart_rx_item_pkg::*;
    import uart_rx_agent_pkg::*;
    import uart_rx_tb_pkg::*;
    

    `include "uart_rx_base_seq.svh"  
           
    `include "uart_rx_input_seq.svh"
   

endpackage : uart_rx_seq_pkg
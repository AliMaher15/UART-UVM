package uart_tx_global_params_pkg;

    parameter DATA_WIDTH = `uart_data_width;
    parameter CLK_PERIOD = `uart_clk_period;
    
endpackage: uart_tx_global_params_pkg
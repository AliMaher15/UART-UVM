package uart_tx_test_pkg ;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import uart_tx_item_pkg::*;
    import uart_tx_global_params_pkg::*;
    import uart_tx_usertypes_pkg::*;
    import uart_tx_agent_pkg::*;
    import uart_tx_seq_pkg::*;
    import uart_tx_tb_pkg::*;

    `include "uart_tx_vseq_base.svh"    
    `include "uart_tx_base_test.svh"

    `include "uart_tx_input_test_vseq.svh"
    `include "uart_tx_input_test.svh"

    `include "active_reset_test.svh"
    `include "idle_reset_test.svh"
    `include "state_transition_reset_test.svh"

endpackage : uart_tx_test_pkg
interface uart_tx_system_if (input clk);

    bit    res_n;    //output
    
endinterface : uart_tx_system_if
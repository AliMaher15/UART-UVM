package uart_tx_global_params_pkg;

    parameter DATA_WIDTH = 8;
    
endpackage: uart_tx_global_params_pkg
package uart_tx_seq_pkg ;
    
	import uvm_pkg::*;
	`include "uvm_macros.svh"

    import uart_tx_item_pkg::*;
    import uart_tx_agent_pkg::*;
    import uart_tx_tb_pkg::*;
    

    `include "uart_tx_base_seq.svh"  
           
    `include "uart_tx_input_seq.svh"
    `include "uart_tx_input_constr_seq.svh"
   

endpackage : uart_tx_seq_pkg
package uart_tx_global_params_pkg;

    parameter DATA_WIDTH = `def_uart_DATA_WIDTH;
    
endpackage: uart_tx_global_params_pkg
package uart_rx_item_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import uart_rx_global_params_pkg::DATA_WIDTH;

    
    `include "uart_rx_item.svh"
  
endpackage : uart_rx_item_pkg
package uart_tx_item_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"
    import uart_tx_global_params_pkg::DATA_WIDTH;
    
    `include "uart_tx_item.svh"
  
endpackage : uart_tx_item_pkg
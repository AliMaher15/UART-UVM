package uart_tx_item_pkg;
    
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    
    `include "uart_tx_item.svh"
  
endpackage : uart_tx_item_pkg
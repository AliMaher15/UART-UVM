interface uart_top_system_if (input clk);

    bit    res_n;    //output
    
endinterface : uart_top_system_if